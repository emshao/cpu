module register66(clk, in_en, in_data, out_data, reset);

    input clk, in_en, reset;
    input [65:0] in_data;
    output [65:0] out_data;

    // wire yesWrite;

    // and whenToWrite(yesWrite, 1'b1, in_en);

    dffe_ref dff0(.q(out_data[0]), .d(in_data[0]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff1(.q(out_data[1]), .d(in_data[1]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff2(.q(out_data[2]), .d(in_data[2]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff3(.q(out_data[3]), .d(in_data[3]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff4(.q(out_data[4]), .d(in_data[4]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff5(.q(out_data[5]), .d(in_data[5]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff6(.q(out_data[6]), .d(in_data[6]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff7(.q(out_data[7]), .d(in_data[7]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff8(.q(out_data[8]), .d(in_data[8]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff9(.q(out_data[9]), .d(in_data[9]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff10(.q(out_data[10]), .d(in_data[10]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff11(.q(out_data[11]), .d(in_data[11]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff12(.q(out_data[12]), .d(in_data[12]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff13(.q(out_data[13]), .d(in_data[13]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff14(.q(out_data[14]), .d(in_data[14]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff15(.q(out_data[15]), .d(in_data[15]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff16(.q(out_data[16]), .d(in_data[16]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff17(.q(out_data[17]), .d(in_data[17]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff18(.q(out_data[18]), .d(in_data[18]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff19(.q(out_data[19]), .d(in_data[19]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff20(.q(out_data[20]), .d(in_data[20]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff21(.q(out_data[21]), .d(in_data[21]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff22(.q(out_data[22]), .d(in_data[22]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff23(.q(out_data[23]), .d(in_data[23]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff24(.q(out_data[24]), .d(in_data[24]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff25(.q(out_data[25]), .d(in_data[25]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff26(.q(out_data[26]), .d(in_data[26]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff27(.q(out_data[27]), .d(in_data[27]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff28(.q(out_data[28]), .d(in_data[28]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff29(.q(out_data[29]), .d(in_data[29]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff30(.q(out_data[30]), .d(in_data[30]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff31(.q(out_data[31]), .d(in_data[31]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff32(.q(out_data[32]), .d(in_data[32]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff33(.q(out_data[33]), .d(in_data[33]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff34(.q(out_data[34]), .d(in_data[34]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff35(.q(out_data[35]), .d(in_data[35]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff36(.q(out_data[36]), .d(in_data[36]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff37(.q(out_data[37]), .d(in_data[37]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff38(.q(out_data[38]), .d(in_data[38]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff39(.q(out_data[39]), .d(in_data[39]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff40(.q(out_data[40]), .d(in_data[40]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff41(.q(out_data[41]), .d(in_data[41]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff42(.q(out_data[42]), .d(in_data[42]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff43(.q(out_data[43]), .d(in_data[43]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff44(.q(out_data[44]), .d(in_data[44]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff45(.q(out_data[45]), .d(in_data[45]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff46(.q(out_data[46]), .d(in_data[46]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff47(.q(out_data[47]), .d(in_data[47]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff48(.q(out_data[48]), .d(in_data[48]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff49(.q(out_data[49]), .d(in_data[49]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff50(.q(out_data[50]), .d(in_data[50]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff51(.q(out_data[51]), .d(in_data[51]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff52(.q(out_data[52]), .d(in_data[52]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff53(.q(out_data[53]), .d(in_data[53]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff54(.q(out_data[54]), .d(in_data[54]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff55(.q(out_data[55]), .d(in_data[55]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff56(.q(out_data[56]), .d(in_data[56]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff57(.q(out_data[57]), .d(in_data[57]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff58(.q(out_data[58]), .d(in_data[58]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff59(.q(out_data[59]), .d(in_data[59]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff60(.q(out_data[60]), .d(in_data[60]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff61(.q(out_data[61]), .d(in_data[61]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff62(.q(out_data[62]), .d(in_data[62]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff63(.q(out_data[63]), .d(in_data[63]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff64(.q(out_data[64]), .d(in_data[64]), .clk(clk), .en(in_en), .clr(reset));
    dffe_ref dff65(.q(out_data[65]), .d(in_data[65]), .clk(clk), .en(in_en), .clr(reset));

    // should be in loop
    // dffe_ref dff0(.q(out_data[0]), .d(in_data[0]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff1(.q(out_data[1]), .d(in_data[1]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff2(.q(out_data[2]), .d(in_data[2]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff3(.q(out_data[3]), .d(in_data[3]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff4(.q(out_data[4]), .d(in_data[4]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff5(.q(out_data[5]), .d(in_data[5]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff6(.q(out_data[6]), .d(in_data[6]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff7(.q(out_data[7]), .d(in_data[7]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff8(.q(out_data[8]), .d(in_data[8]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff9(.q(out_data[9]), .d(in_data[9]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff10(.q(out_data[10]), .d(in_data[10]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff11(.q(out_data[11]), .d(in_data[11]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff12(.q(out_data[12]), .d(in_data[12]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff13(.q(out_data[13]), .d(in_data[13]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff14(.q(out_data[14]), .d(in_data[14]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff15(.q(out_data[15]), .d(in_data[15]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff16(.q(out_data[16]), .d(in_data[16]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff17(.q(out_data[17]), .d(in_data[17]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff18(.q(out_data[18]), .d(in_data[18]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff19(.q(out_data[19]), .d(in_data[19]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff20(.q(out_data[20]), .d(in_data[20]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff21(.q(out_data[21]), .d(in_data[21]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff22(.q(out_data[22]), .d(in_data[22]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff23(.q(out_data[23]), .d(in_data[23]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff24(.q(out_data[24]), .d(in_data[24]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff25(.q(out_data[25]), .d(in_data[25]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff26(.q(out_data[26]), .d(in_data[26]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff27(.q(out_data[27]), .d(in_data[27]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff28(.q(out_data[28]), .d(in_data[28]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff29(.q(out_data[29]), .d(in_data[29]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff30(.q(out_data[30]), .d(in_data[30]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff31(.q(out_data[31]), .d(in_data[31]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff32(.q(out_data[32]), .d(in_data[32]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff33(.q(out_data[33]), .d(in_data[33]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff34(.q(out_data[34]), .d(in_data[34]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff35(.q(out_data[35]), .d(in_data[35]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff36(.q(out_data[36]), .d(in_data[36]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff37(.q(out_data[37]), .d(in_data[37]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff38(.q(out_data[38]), .d(in_data[38]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff39(.q(out_data[39]), .d(in_data[39]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff40(.q(out_data[40]), .d(in_data[40]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff41(.q(out_data[41]), .d(in_data[41]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff42(.q(out_data[42]), .d(in_data[42]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff43(.q(out_data[43]), .d(in_data[43]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff44(.q(out_data[44]), .d(in_data[44]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff45(.q(out_data[45]), .d(in_data[45]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff46(.q(out_data[46]), .d(in_data[46]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff47(.q(out_data[47]), .d(in_data[47]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff48(.q(out_data[48]), .d(in_data[48]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff49(.q(out_data[49]), .d(in_data[49]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff50(.q(out_data[50]), .d(in_data[50]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff51(.q(out_data[51]), .d(in_data[51]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff52(.q(out_data[52]), .d(in_data[52]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff53(.q(out_data[53]), .d(in_data[53]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff54(.q(out_data[54]), .d(in_data[54]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff55(.q(out_data[55]), .d(in_data[55]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff56(.q(out_data[56]), .d(in_data[56]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff57(.q(out_data[57]), .d(in_data[57]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff58(.q(out_data[58]), .d(in_data[58]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff59(.q(out_data[59]), .d(in_data[59]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff60(.q(out_data[60]), .d(in_data[60]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff61(.q(out_data[61]), .d(in_data[61]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff62(.q(out_data[62]), .d(in_data[62]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff63(.q(out_data[63]), .d(in_data[63]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff64(.q(out_data[64]), .d(in_data[64]), .clk(clk), .en(yesWrite), .clr(reset));
    // dffe_ref dff65(.q(out_data[65]), .d(in_data[65]), .clk(clk), .en(yesWrite), .clr(reset));


endmodule